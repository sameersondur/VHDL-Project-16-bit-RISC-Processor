library ieee;
use ieee.std_logic_1164.all;

---------Package Declaration-----------------------------------
package arr is 
  type array_rom is array (0 to 255) of std_logic_vector(15 downto 0); -- subtype for ROM
end package arr;
----------------------------------------------------------------


use  work.arr.all;
library ieee;
use ieee.std_logic_1164.all;
USE ieee.numeric_std.ALL;

--------------Entity Declaration ---------------------
entity instruction_memory is 
  port( pc: in std_logic_vector(7 downto 0);
        instruction: out std_logic_vector(15 downto 0));  
end entity instruction_memory;
-------------------------------------------------------

-------------Architecture Body Declaration------------------
architecture arch_instr_mem of instruction_memory is
  signal ROM: array_rom;
begin  
ROM(0) <=   "0001000000001111" ; -- ADD R[0], #00001111
ROM(1) <=   "0111000100000010";	-- interrupt enable
ROM(2) <=   "0010000000000001";  -- ADD R[0], R[1]
ROM(3) <=   "0100000000000001"; -- SHL R[0], R[1]
ROM(4) <=   "0001001010101010"; -- ADD R[2], #10101010
ROM(5) <=   "0001001110101010"; -- ADD R[3], #10101010
ROM(6) <=   "0101001100100011"; -- XOR R[2], R[3]
ROM(7) <=   "1000000001000000"; -- LD R[4], Mem[0]
ROM(8) <=   "0001111100000001"; -- immed R[15],0001
ROM(9) <=   "0001010000001001"; -- immed R[4], 1001
ROM(10) <=  "1001000000010100"; -- STR Mem[1], R[4]
ROM(11) <=  "1000000001010001"; -- LD R[5], mem[1]
ROM(12) <=  "0010000001010010"; -- Add R[5],R[2]  check value of rx from earlier thing
ROM(13) <=  "0101011000010000"; -- CLR R[1]
ROM(14) <=  "0101010100010010"; -- OR R[1], R[2]
ROM(15) <=  "0101100000010010"; -- MOV R[1], R[2]
ROM(16) <=  "0101011000110000"; -- CLR R[3]
ROM(17) <=  "1101000000110100"; -- JZ #0100
ROM(18) <=   "0000000000000000"; -- NOP
ROM(19) <=  "0101011101000000"; -- SET R[4]
ROM(20) <=  "1110000001000001"; -- JNZ #0001
ROM(21) <=   "0000000000000000"; -- NOP
ROM(22) <=   "1010000000000001"; -- LD R[0], #0001
ROM(23) <=   "1011000100000010"; -- STR #0010 , R[1]
ROM(24) <=  "0101011101100000"; -- SET R[6]
ROM(25) <=   "0001011100000001"; -- ADD R[7], 00000001
ROM(26) <=   "0001100000000100"; -- ADD R[8], 00000100
ROM(27) <=   "0101111101111000"; -- SLT R[7], R[8]
ROM(28) <=   "0011000101110000"; -- DEC R[7]
ROM(29) <=  "0101000001110000"; -- NOT R[7]
ROM(30) <=  "0101000101111000"; -- NOR R[7], R[8]
ROM(31) <=  "0101010001111000" ; -- AND R[7], R[8]
ROM(32) <=   "1100000000000001"; -- JMP #00000001

ROM(128)<="0001000000001111" ; -- ADD R[0], #00001111
ROM(129)<="0001000100000010";	-- ADD R[1], #00000010
ROM(130)<= "0010000000000001";  -- ADD R[0], R[1]
ROM(131) <=   "0100000000000001"; -- SHL R[0], R[1]
ROM(132) <=   "0001001010101010"; -- ADD R[2], #10101010
ROM(133) <=   "0001001110101010"; -- ADD R[3], #10101010
ROM(134) <=   "1111000001000000"; -- return
ROM(135) <=   "0000000000000000"; -- return

ROM(153)<="0001000000001111" ; -- ADD R[0], #00001111
ROM(154)<="0001000100000010";	-- ADD R[1], #00000010
ROM(155)<= "0010000000000001";  -- ADD R[0], R[1]
ROM(156) <=   "0100000000000001"; -- SHL R[0], R[1]
ROM(157) <=   "0001001010101010"; -- ADD R[2], #10101010
ROM(158) <=   "0001001110101010"; -- ADD R[3], #10101010
ROM(159) <=   "1111000001000000"; -- return
ROM(160) <=   "0000000000000000"; -- return

ROM(178)<="0001111100001111" ; -- ADD R[15], #00001111
ROM(179)<="0001101000000010";	-- ADD R[10], #00000010
ROM(180)<= "0010000010101111";  -- ADD R[10], R[15]
ROM(181) <= "0101000001110000"; -- NOT R[7]
ROM(182) <=   "0001010110101010"; -- ADD R[5], #10101010
ROM(183) <=   "1111000001000000"; -- return
ROM(184) <=   "0000000000000000"; -- return

ROM(203)<="0101011101000000"; -- SET R[4]
ROM(204)<="0001010000000010";	-- ADD R[4], #00000010
ROM(205)<= "0010000010101111";  -- ADD R[10], R[15]
ROM(206) <= "0101000001110000"; -- NOT R[7]
ROM(207) <=  "0101010001111000" ; -- AND R[7], R[8]
ROM(208) <=   "1111000001000000"; -- return
ROM(209) <=   "0000000000000000"; -- return

  --------Process Declaration----------------------
  seq: process (pc) is
  begin
    instruction <= ROM (to_integer(unsigned(pc)));     
 end process seq;
 ----------------------------------------------------
 
end architecture arch_instr_mem;    --architecture ends here
